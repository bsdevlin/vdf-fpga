/*
  Copyright (C) 2019  Benjamin Devlin

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
 */

/*
 This performs repeated modular squaring using Montgomery multiplication technique.

 We use redundant bit representation to minimize delay from carry chains.

 Single clock cycle multiplier which can either calculate the square, lower, or upper
 products is used.

 Montgomery parameters are extended to include a redundant word so that we can skip the final
 overflow check.

 One hot control signals.

 Everything fits inside a single SLR.

 redun_mont_pkg contains functions for calculating Montgomery values and commonly used typedefs.
 */

module redun_mont
  import redun_mont_pkg::*;
(
  input           i_clk,
  input           i_rst,
  input redun0_t  i_sq,
  input           i_val,
  output redun0_t o_mul,
  output logic    o_val
);

redun0_t mul_a, mul_b, hmul_out_h, hmul_out_h_r, tmp_h, i_sq_r, i_sq_rr, mult_out_l, mult_out_l_r;
redun1_t mult_out, mult_out_r;

logic [63:0] ovrflw_cnt;
logic o_val_r, i_val_r;

typedef enum logic [5:0] {IDLE  = 1 << 0,
                          START = 1 << 1,
                          MUL0  = 2 << 1,
                          MUL1  = 3 << 1,
                          MUL2  = 4 << 1,
                          MUL2_OVRFLW = 5 << 1} state_index_t;
                          
state_index_t state, state_r, next_state;
      
typedef enum logic [2:0] {SQR  = 1 << 0,
                          MUL_L = 1 << 1,
                          MUL_H  = 1 << 2} mult_ctl_t;     
      
mult_ctl_t mult_ctl, next_mult_ctl; 


// Assign input to multiplier
always_comb begin
  for (int i = 0; i < NUM_WRDS; i++)
    hmul_out_h[i] = mult_out[NUM_WRDS-1-i];

  mult_out_l = mult_out[0:NUM_WRDS-1];

  mul_a = i_sq_rr;
  mul_b = i_sq_rr;

  unique case (state)
    IDLE: begin
      mul_a = i_sq_rr;
      mul_b = i_sq_rr;
      next_mult_ctl = SQR;
      if (i_val_r)
        next_state = START;
      else
        next_state = IDLE;
    end
    START: begin
      mul_a = i_sq_rr;
      mul_b = i_sq_rr;
      next_state = MUL0;
      next_mult_ctl = MUL_L;
    end
    MUL0: begin
      mul_a = mult_out_l;
      mul_b = to_redun(MONT_FACTOR);
      next_mult_ctl = MUL_H;
      if (&mult_out[NUM_WRDS][WRD_BITS-1:0])
        next_state = MUL2_OVRFLW;
      else
        next_state = MUL1;
    end
    MUL1: begin
      mul_a = mult_out_l;
      mul_a[NUM_WRDS-1][WRD_BITS] = 0; // what if we had 0xffff - TODO
      mul_b = to_redun(P);
      next_state = MUL2;
      next_mult_ctl = SQR;
    end
    MUL2: begin
      mul_a = hmul_out_h;
      mul_b = hmul_out_h;
      
      next_state = MUL0;
      next_mult_ctl = MUL_L;
      
      // Need to do low multiplication if we detect possible overflow
      if (&mult_out[NUM_WRDS][WRD_BITS-1:0]) begin
        next_state = MUL2_OVRFLW;
        next_mult_ctl = MUL_L;
      end
    end
    // Here we calculate the lower words to check for overflow
    MUL2_OVRFLW: begin
      mul_a = mult_out_l_r;
      mul_a[NUM_WRDS-1][WRD_BITS] = 0;
      mul_b = to_redun(P);
      next_mult_ctl = MUL_L;
      next_state = MUL2_OVRFLW;
      if (state_r == MUL2_OVRFLW && ~(&mult_out[NUM_WRDS-2][WRD_BITS-1:0])) begin
        next_state = START;
        next_mult_ctl = SQR;
      end
    end
  endcase
end

// Logic without a reset
always_ff @ (posedge i_clk) begin
  state_r <= state;
  i_sq_r <= i_sq;
  if (state == MUL0)
    for (int i = 0; i < NUM_WRDS; i++)
      tmp_h[i] <= mult_out[NUM_WRDS+i] + (i == 0 ? (mult_out[NUM_WRDS-1][WRD_BITS] + 1) : 0);
  else
    tmp_h <= to_redun(0);
  
  mult_ctl <= next_mult_ctl;
  mult_out_r <= mult_out;
  if (state == MUL1)
    mult_out_l_r <= mult_out_l;
    
  i_val_r <= i_val;
  o_val_r <= state == MUL2 && state_r != MUL2_OVRFLW;
  o_val <= o_val_r;
      
  // Here we do the overflow check for mul2
  if (state == MUL2_OVRFLW) begin
    o_val_r <= next_state != MUL2_OVRFLW;
    
    o_val <= 0;
    if (state_r == MUL2_OVRFLW)
      for (int i = 0; i < NUM_WRDS; i++) begin
        i_sq_rr[i] <= i_sq_rr[i][WRD_BITS-1:0] + (i == 0 ? mult_out[NUM_WRDS-2][WRD_BITS] : i_sq_rr[i-1][WRD_BITS]);
        hmul_out_h_r[i] <= hmul_out_h_r[i][WRD_BITS-1:0] + (i == 0 ? mult_out[NUM_WRDS-2][WRD_BITS] : hmul_out_h_r[i-1][WRD_BITS]);
      end
  end else begin
    i_sq_rr <= hmul_out_h;
    hmul_out_h_r <= hmul_out_h;
    o_mul <= hmul_out_h_r;
  end
  
  if (state == IDLE)
    i_sq_rr <= i_sq_r;

end

// Logic requiring reset
always_ff @ (posedge i_clk) begin
  if (i_rst) begin
    state <= IDLE;
    ovrflw_cnt <= 0;
  end else begin
    state <= next_state;
    if (state == MUL2_OVRFLW && state_r != MUL2_OVRFLW)
      ovrflw_cnt <= ovrflw_cnt + 1;
  end
end

multi_mode_multiplier #(
  .NUM_ELEMENTS    ( NUM_WRDS                        ),
  .DSP_BIT_LEN     ( WRD_BITS+1                      ),
  .WORD_LEN        ( WRD_BITS                        ),
  .NUM_ELEMENTS_OUT( NUM_WRDS+SPECULATIVE_CARRY_WRDS )
)
multi_mode_multiplier (
  .i_clk      ( i_clk    ),
  .i_ctl      ( mult_ctl ),
  .i_dat_a    ( mul_a    ),
  .i_dat_b    ( mul_b    ),
  .i_add_term ( tmp_h    ),
  .o_dat      ( mult_out )
);

endmodule
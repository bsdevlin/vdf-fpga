
// Coef 0
always_ff @ (posedge i_clk) accum_grid_o[0] <= {{1{1'd0}},mul_grid[0][0][0+:17],{0{1'd0}}};

// Coef 1
logic [18:0] accum_i_1 [3];
logic [18:0] accum_o_c_1, accum_o_s_1;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(3),
  .BIT_LEN(19)
)
ct_1 (
  .terms(accum_i_1),
  .C(accum_o_c_1),
  .S(accum_o_s_1)
);
always_comb accum_i_1 = {{{0{1'd0}},mul_grid[0][0][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][1][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][0][0+:8],{9{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[1] <= accum_o_c_1 + accum_o_s_1;

// Coef 2
logic [19:0] accum_i_2 [5];
logic [19:0] accum_o_c_2, accum_o_s_2;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(5),
  .BIT_LEN(20)
)
ct_2 (
  .terms(accum_i_2),
  .C(accum_o_c_2),
  .S(accum_o_s_2)
);
always_comb accum_i_2 = {{{0{1'd0}},mul_grid[0][0][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][1][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][2][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][0][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][1][0+:8],{9{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[2] <= accum_o_c_2 + accum_o_s_2;

// Coef 3
logic [19:0] accum_i_3 [7];
logic [19:0] accum_o_c_3, accum_o_s_3;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(7),
  .BIT_LEN(20)
)
ct_3 (
  .terms(accum_i_3),
  .C(accum_o_c_3),
  .S(accum_o_s_3)
);
always_comb accum_i_3 = {{{0{1'd0}},mul_grid[0][1][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][2][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][3][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][0][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][1][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][2][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][0][0+:16],{1{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[3] <= accum_o_c_3 + accum_o_s_3;

// Coef 4
logic [20:0] accum_i_4 [10];
logic [20:0] accum_o_c_4, accum_o_s_4;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(10),
  .BIT_LEN(21)
)
ct_4 (
  .terms(accum_i_4),
  .C(accum_o_c_4),
  .S(accum_o_s_4)
);
always_comb accum_i_4 = {{{0{1'd0}},mul_grid[0][2][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][3][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][4][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][0][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][1][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][2][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][3][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][0][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][1][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][0][0+:7],{10{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[4] <= accum_o_c_4 + accum_o_s_4;

// Coef 5
logic [20:0] accum_i_5 [12];
logic [20:0] accum_o_c_5, accum_o_s_5;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(12),
  .BIT_LEN(21)
)
ct_5 (
  .terms(accum_i_5),
  .C(accum_o_c_5),
  .S(accum_o_s_5)
);
always_comb accum_i_5 = {{{0{1'd0}},mul_grid[0][3][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][4][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][5][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][1][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][2][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][3][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][4][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][0][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][1][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][2][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][0][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][1][0+:7],{10{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[5] <= accum_o_c_5 + accum_o_s_5;

// Coef 6
logic [20:0] accum_i_6 [14];
logic [20:0] accum_o_c_6, accum_o_s_6;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(14),
  .BIT_LEN(21)
)
ct_6 (
  .terms(accum_i_6),
  .C(accum_o_c_6),
  .S(accum_o_s_6)
);
always_comb accum_i_6 = {{{0{1'd0}},mul_grid[0][4][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][5][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][6][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][2][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][3][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][4][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][5][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][1][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][2][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][3][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][0][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][1][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][2][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][0][0+:15],{2{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[6] <= accum_o_c_6 + accum_o_s_6;

// Coef 7
logic [20:0] accum_i_7 [17];
logic [20:0] accum_o_c_7, accum_o_s_7;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(17),
  .BIT_LEN(21)
)
ct_7 (
  .terms(accum_i_7),
  .C(accum_o_c_7),
  .S(accum_o_s_7)
);
always_comb accum_i_7 = {{{0{1'd0}},mul_grid[0][5][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][6][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][7][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][3][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][4][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][5][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][6][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][2][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][3][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][4][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][0][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][1][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][2][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][3][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][0][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][1][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][0][0+:6],{11{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[7] <= accum_o_c_7 + accum_o_s_7;

// Coef 8
logic [21:0] accum_i_8 [19];
logic [21:0] accum_o_c_8, accum_o_s_8;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(19),
  .BIT_LEN(22)
)
ct_8 (
  .terms(accum_i_8),
  .C(accum_o_c_8),
  .S(accum_o_s_8)
);
always_comb accum_i_8 = {{{0{1'd0}},mul_grid[0][6][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][7][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][8][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][4][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][5][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][6][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][7][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][3][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][4][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][5][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][1][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][2][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][3][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][4][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][0][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][1][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][2][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][0][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][1][0+:6],{11{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[8] <= accum_o_c_8 + accum_o_s_8;

// Coef 9
logic [21:0] accum_i_9 [21];
logic [21:0] accum_o_c_9, accum_o_s_9;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(21),
  .BIT_LEN(22)
)
ct_9 (
  .terms(accum_i_9),
  .C(accum_o_c_9),
  .S(accum_o_s_9)
);
always_comb accum_i_9 = {{{0{1'd0}},mul_grid[0][7][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][8][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][9][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][5][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][6][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][7][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][8][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][4][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][5][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][6][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][2][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][3][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][4][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][5][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][1][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][2][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][3][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][0][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][1][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][2][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][0][0+:14],{3{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[9] <= accum_o_c_9 + accum_o_s_9;

// Coef 10
logic [21:0] accum_i_10 [24];
logic [21:0] accum_o_c_10, accum_o_s_10;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(24),
  .BIT_LEN(22)
)
ct_10 (
  .terms(accum_i_10),
  .C(accum_o_c_10),
  .S(accum_o_s_10)
);
always_comb accum_i_10 = {{{0{1'd0}},mul_grid[0][8][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][9][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][10][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][6][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][7][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][8][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][9][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][5][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][6][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][7][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][3][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][4][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][5][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][6][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][2][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][3][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][4][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][0][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][1][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][2][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][3][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][0][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][1][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][0][0+:5],{12{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[10] <= accum_o_c_10 + accum_o_s_10;

// Coef 11
logic [21:0] accum_i_11 [26];
logic [21:0] accum_o_c_11, accum_o_s_11;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(26),
  .BIT_LEN(22)
)
ct_11 (
  .terms(accum_i_11),
  .C(accum_o_c_11),
  .S(accum_o_s_11)
);
always_comb accum_i_11 = {{{0{1'd0}},mul_grid[0][9][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][10][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][11][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][7][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][8][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][9][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][10][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][6][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][7][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][8][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][4][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][5][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][6][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][7][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][3][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][4][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][5][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][1][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][2][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][3][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][4][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][0][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][1][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][2][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][0][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][1][0+:5],{12{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[11] <= accum_o_c_11 + accum_o_s_11;

// Coef 12
logic [21:0] accum_i_12 [28];
logic [21:0] accum_o_c_12, accum_o_s_12;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(28),
  .BIT_LEN(22)
)
ct_12 (
  .terms(accum_i_12),
  .C(accum_o_c_12),
  .S(accum_o_s_12)
);
always_comb accum_i_12 = {{{0{1'd0}},mul_grid[0][10][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][11][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][12][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][8][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][9][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][10][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][11][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][7][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][8][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][9][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][5][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][6][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][7][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][8][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][4][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][5][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][6][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][2][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][3][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][4][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][5][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][1][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][2][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][3][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][0][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][1][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][2][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][0][0+:13],{4{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[12] <= accum_o_c_12 + accum_o_s_12;

// Coef 13
logic [21:0] accum_i_13 [31];
logic [21:0] accum_o_c_13, accum_o_s_13;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(31),
  .BIT_LEN(22)
)
ct_13 (
  .terms(accum_i_13),
  .C(accum_o_c_13),
  .S(accum_o_s_13)
);
always_comb accum_i_13 = {{{0{1'd0}},mul_grid[0][11][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][12][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][13][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][9][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][10][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][11][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][12][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][8][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][9][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][10][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][6][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][7][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][8][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][9][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][5][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][6][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][7][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][3][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][4][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][5][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][6][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][2][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][3][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][4][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][0][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][1][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][2][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][3][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][0][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][1][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][0][0+:4],{13{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[13] <= accum_o_c_13 + accum_o_s_13;

// Coef 14
logic [21:0] accum_i_14 [33];
logic [21:0] accum_o_c_14, accum_o_s_14;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(33),
  .BIT_LEN(22)
)
ct_14 (
  .terms(accum_i_14),
  .C(accum_o_c_14),
  .S(accum_o_s_14)
);
always_comb accum_i_14 = {{{0{1'd0}},mul_grid[0][12][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][13][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][14][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][10][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][11][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][12][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][13][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][9][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][10][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][11][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][7][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][8][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][9][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][10][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][6][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][7][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][8][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][4][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][5][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][6][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][7][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][3][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][4][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][5][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][1][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][2][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][3][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][4][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][0][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][1][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][2][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][0][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][1][0+:4],{13{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[14] <= accum_o_c_14 + accum_o_s_14;

// Coef 15
logic [21:0] accum_i_15 [35];
logic [21:0] accum_o_c_15, accum_o_s_15;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(35),
  .BIT_LEN(22)
)
ct_15 (
  .terms(accum_i_15),
  .C(accum_o_c_15),
  .S(accum_o_s_15)
);
always_comb accum_i_15 = {{{0{1'd0}},mul_grid[0][13][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][14][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][15][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][11][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][12][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][13][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][14][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][10][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][11][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][12][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][8][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][9][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][10][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][11][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][7][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][8][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][9][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][5][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][6][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][7][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][8][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][4][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][5][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][6][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][2][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][3][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][4][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][5][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][1][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][2][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][3][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][0][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][1][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][2][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][0][0+:12],{5{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[15] <= accum_o_c_15 + accum_o_s_15;

// Coef 16
logic [22:0] accum_i_16 [38];
logic [22:0] accum_o_c_16, accum_o_s_16;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(38),
  .BIT_LEN(23)
)
ct_16 (
  .terms(accum_i_16),
  .C(accum_o_c_16),
  .S(accum_o_s_16)
);
always_comb accum_i_16 = {{{0{1'd0}},mul_grid[0][14][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][15][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][16][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][12][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][13][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][14][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][15][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][11][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][12][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][13][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][9][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][10][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][11][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][12][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][8][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][9][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][10][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][6][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][7][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][8][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][9][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][5][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][6][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][7][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][3][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][4][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][5][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][6][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][2][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][3][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][4][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][0][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][1][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][2][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][3][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][0][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][1][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][0][0+:3],{14{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[16] <= accum_o_c_16 + accum_o_s_16;

// Coef 17
logic [22:0] accum_i_17 [40];
logic [22:0] accum_o_c_17, accum_o_s_17;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(40),
  .BIT_LEN(23)
)
ct_17 (
  .terms(accum_i_17),
  .C(accum_o_c_17),
  .S(accum_o_s_17)
);
always_comb accum_i_17 = {{{0{1'd0}},mul_grid[0][15][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][16][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][17][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][13][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][14][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][15][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][16][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][12][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][13][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][14][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][10][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][11][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][12][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][13][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][9][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][10][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][11][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][7][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][8][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][9][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][10][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][6][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][7][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][8][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][4][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][5][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][6][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][7][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][3][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][4][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][5][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][1][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][2][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][3][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][4][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][0][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][1][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][2][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][0][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][1][0+:3],{14{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[17] <= accum_o_c_17 + accum_o_s_17;

// Coef 18
logic [22:0] accum_i_18 [42];
logic [22:0] accum_o_c_18, accum_o_s_18;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(42),
  .BIT_LEN(23)
)
ct_18 (
  .terms(accum_i_18),
  .C(accum_o_c_18),
  .S(accum_o_s_18)
);
always_comb accum_i_18 = {{{0{1'd0}},mul_grid[0][16][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][17][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][18][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][14][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][15][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][16][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][17][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][13][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][14][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][15][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][11][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][12][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][13][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][14][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][10][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][11][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][12][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][8][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][9][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][10][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][11][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][7][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][8][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][9][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][5][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][6][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][7][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][8][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][4][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][5][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][6][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][2][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][3][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][4][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][5][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][1][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][2][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][3][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][0][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][1][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][2][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][0][0+:11],{6{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[18] <= accum_o_c_18 + accum_o_s_18;

// Coef 19
logic [22:0] accum_i_19 [45];
logic [22:0] accum_o_c_19, accum_o_s_19;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(45),
  .BIT_LEN(23)
)
ct_19 (
  .terms(accum_i_19),
  .C(accum_o_c_19),
  .S(accum_o_s_19)
);
always_comb accum_i_19 = {{{0{1'd0}},mul_grid[0][17][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][18][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][19][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][15][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][16][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][17][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][18][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][14][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][15][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][16][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][12][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][13][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][14][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][15][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][11][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][12][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][13][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][9][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][10][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][11][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][12][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][8][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][9][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][10][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][6][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][7][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][8][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][9][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][5][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][6][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][7][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][3][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][4][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][5][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][6][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][2][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][3][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][4][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][0][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][1][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][2][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][3][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][0][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][1][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][0][0+:2],{15{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[19] <= accum_o_c_19 + accum_o_s_19;

// Coef 20
logic [22:0] accum_i_20 [47];
logic [22:0] accum_o_c_20, accum_o_s_20;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(47),
  .BIT_LEN(23)
)
ct_20 (
  .terms(accum_i_20),
  .C(accum_o_c_20),
  .S(accum_o_s_20)
);
always_comb accum_i_20 = {{{0{1'd0}},mul_grid[0][18][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][19][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][20][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][16][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][17][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][18][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][19][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][15][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][16][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][17][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][13][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][14][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][15][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][16][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][12][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][13][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][14][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][10][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][11][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][12][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][13][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][9][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][10][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][11][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][7][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][8][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][9][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][10][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][6][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][7][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][8][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][4][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][5][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][6][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][7][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][3][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][4][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][5][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][1][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][2][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][3][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][4][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][0][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][1][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][2][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][0][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][1][0+:2],{15{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[20] <= accum_o_c_20 + accum_o_s_20;

// Coef 21
logic [22:0] accum_i_21 [49];
logic [22:0] accum_o_c_21, accum_o_s_21;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(49),
  .BIT_LEN(23)
)
ct_21 (
  .terms(accum_i_21),
  .C(accum_o_c_21),
  .S(accum_o_s_21)
);
always_comb accum_i_21 = {{{0{1'd0}},mul_grid[0][19][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][20][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][21][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][17][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][18][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][19][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][20][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][16][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][17][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][18][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][14][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][15][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][16][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][17][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][13][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][14][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][15][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][11][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][12][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][13][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][14][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][10][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][11][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][12][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][8][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][9][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][10][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][11][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][7][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][8][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][9][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][5][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][6][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][7][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][8][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][4][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][5][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][6][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][2][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][3][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][4][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][5][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][1][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][2][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][3][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][0][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][1][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][2][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][0][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[21] <= accum_o_c_21 + accum_o_s_21;

// Coef 22
logic [22:0] accum_i_22 [51];
logic [22:0] accum_o_c_22, accum_o_s_22;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(51),
  .BIT_LEN(23)
)
ct_22 (
  .terms(accum_i_22),
  .C(accum_o_c_22),
  .S(accum_o_s_22)
);
always_comb accum_i_22 = {{{0{1'd0}},mul_grid[0][20][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][21][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[0][22][0+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][18][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][19][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][20][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][21][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][17][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][18][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][19][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][15][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][16][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][17][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][18][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][14][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][15][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][16][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][12][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][13][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][14][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][15][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][11][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][12][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][13][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][9][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][10][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][11][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][12][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][8][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][9][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][10][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][6][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][7][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][8][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][9][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][5][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][6][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][7][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][3][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][4][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][5][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][6][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][2][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][3][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][4][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][0][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][1][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][2][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][3][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][0][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][1][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[22] <= accum_o_c_22 + accum_o_s_22;

// Coef 23
logic [22:0] accum_i_23 [51];
logic [22:0] accum_o_c_23, accum_o_s_23;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(51),
  .BIT_LEN(23)
)
ct_23 (
  .terms(accum_i_23),
  .C(accum_o_c_23),
  .S(accum_o_s_23)
);
always_comb accum_i_23 = {{{0{1'd0}},mul_grid[0][21][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[0][22][17+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][19][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][20][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][21][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][22][0+:8],{9{1'd0}}},{{0{1'd0}},mul_grid[2][18][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][19][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][20][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][16][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][17][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][18][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][19][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][15][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][16][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][17][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][13][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][14][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][15][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][16][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][12][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][13][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][14][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][10][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][11][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][12][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][13][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][9][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][10][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][11][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][7][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][8][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][9][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][10][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][6][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][7][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][8][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][4][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][5][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][6][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][7][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][3][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][4][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][5][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][1][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][2][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][3][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][4][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][0][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][1][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][2][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[23] <= accum_o_c_23 + accum_o_s_23;

// Coef 24
logic [22:0] accum_i_24 [49];
logic [22:0] accum_o_c_24, accum_o_s_24;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(49),
  .BIT_LEN(23)
)
ct_24 (
  .terms(accum_i_24),
  .C(accum_o_c_24),
  .S(accum_o_s_24)
);
always_comb accum_i_24 = {{{0{1'd0}},mul_grid[0][22][34+:9],{0{1'd0}}},{{0{1'd0}},mul_grid[1][20][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][21][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[1][22][8+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][19][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][20][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][21][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][17][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][18][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][19][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][20][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][16][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][17][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][18][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][14][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][15][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][16][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][17][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][13][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][14][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][15][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][11][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][12][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][13][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][14][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][10][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][11][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][12][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][8][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][9][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][10][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][11][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][7][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][8][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][9][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][5][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][6][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][7][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][8][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][4][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][5][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][6][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][2][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][3][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][4][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][5][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][1][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][2][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][3][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[24] <= accum_o_c_24 + accum_o_s_24;

// Coef 25
logic [22:0] accum_i_25 [47];
logic [22:0] accum_o_c_25, accum_o_s_25;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(47),
  .BIT_LEN(23)
)
ct_25 (
  .terms(accum_i_25),
  .C(accum_o_c_25),
  .S(accum_o_s_25)
);
always_comb accum_i_25 = {{{0{1'd0}},mul_grid[1][21][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[1][22][25+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][20][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][21][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[2][22][0+:16],{1{1'd0}}},{{0{1'd0}},mul_grid[3][18][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][19][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][20][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][21][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][17][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][18][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][19][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][15][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][16][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][17][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][18][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][14][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][15][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][16][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][12][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][13][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][14][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][15][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][11][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][12][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][13][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][9][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][10][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][11][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][12][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][8][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][9][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][10][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][6][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][7][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][8][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][9][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][5][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][6][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][7][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][3][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][4][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][5][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][6][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][2][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][3][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][4][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[25] <= accum_o_c_25 + accum_o_s_25;

// Coef 26
logic [22:0] accum_i_26 [45];
logic [22:0] accum_o_c_26, accum_o_s_26;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(45),
  .BIT_LEN(23)
)
ct_26 (
  .terms(accum_i_26),
  .C(accum_o_c_26),
  .S(accum_o_s_26)
);
always_comb accum_i_26 = {{{0{1'd0}},mul_grid[1][22][42+:1],{0{1'd0}}},{{0{1'd0}},mul_grid[2][21][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[2][22][16+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][19][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][20][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][21][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][22][0+:7],{10{1'd0}}},{{0{1'd0}},mul_grid[4][18][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][19][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][20][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][16][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][17][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][18][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][19][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][15][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][16][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][17][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][13][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][14][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][15][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][16][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][12][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][13][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][14][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][10][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][11][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][12][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][13][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][9][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][10][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][11][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][7][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][8][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][9][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][10][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][6][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][7][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][8][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][4][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][5][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][6][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][7][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][3][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][4][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][5][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[26] <= accum_o_c_26 + accum_o_s_26;

// Coef 27
logic [22:0] accum_i_27 [42];
logic [22:0] accum_o_c_27, accum_o_s_27;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(42),
  .BIT_LEN(23)
)
ct_27 (
  .terms(accum_i_27),
  .C(accum_o_c_27),
  .S(accum_o_s_27)
);
always_comb accum_i_27 = {{{0{1'd0}},mul_grid[2][22][33+:10],{0{1'd0}}},{{0{1'd0}},mul_grid[3][20][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][21][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[3][22][7+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][19][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][20][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][21][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][17][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][18][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][19][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][20][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][16][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][17][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][18][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][14][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][15][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][16][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][17][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][13][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][14][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][15][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][11][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][12][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][13][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][14][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][10][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][11][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][12][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][8][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][9][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][10][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][11][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][7][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][8][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][9][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][5][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][6][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][7][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][8][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][4][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][5][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][6][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[27] <= accum_o_c_27 + accum_o_s_27;

// Coef 28
logic [22:0] accum_i_28 [40];
logic [22:0] accum_o_c_28, accum_o_s_28;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(40),
  .BIT_LEN(23)
)
ct_28 (
  .terms(accum_i_28),
  .C(accum_o_c_28),
  .S(accum_o_s_28)
);
always_comb accum_i_28 = {{{0{1'd0}},mul_grid[3][21][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[3][22][24+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][20][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][21][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[4][22][0+:15],{2{1'd0}}},{{0{1'd0}},mul_grid[5][18][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][19][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][20][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][21][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][17][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][18][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][19][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][15][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][16][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][17][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][18][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][14][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][15][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][16][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][12][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][13][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][14][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][15][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][11][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][12][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][13][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][9][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][10][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][11][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][12][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][8][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][9][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][10][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][6][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][7][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][8][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][9][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][5][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][6][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][7][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[28] <= accum_o_c_28 + accum_o_s_28;

// Coef 29
logic [21:0] accum_i_29 [38];
logic [21:0] accum_o_c_29, accum_o_s_29;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(38),
  .BIT_LEN(22)
)
ct_29 (
  .terms(accum_i_29),
  .C(accum_o_c_29),
  .S(accum_o_s_29)
);
always_comb accum_i_29 = {{{0{1'd0}},mul_grid[3][22][41+:2],{0{1'd0}}},{{0{1'd0}},mul_grid[4][21][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[4][22][15+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][19][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][20][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][21][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][22][0+:6],{11{1'd0}}},{{0{1'd0}},mul_grid[6][18][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][19][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][20][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][16][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][17][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][18][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][19][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][15][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][16][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][17][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][13][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][14][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][15][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][16][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][12][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][13][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][14][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][10][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][11][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][12][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][13][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][9][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][10][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][11][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][7][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][8][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][9][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][10][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][6][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][7][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][8][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[29] <= accum_o_c_29 + accum_o_s_29;

// Coef 30
logic [21:0] accum_i_30 [35];
logic [21:0] accum_o_c_30, accum_o_s_30;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(35),
  .BIT_LEN(22)
)
ct_30 (
  .terms(accum_i_30),
  .C(accum_o_c_30),
  .S(accum_o_s_30)
);
always_comb accum_i_30 = {{{0{1'd0}},mul_grid[4][22][32+:11],{0{1'd0}}},{{0{1'd0}},mul_grid[5][20][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][21][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[5][22][6+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][19][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][20][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][21][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][17][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][18][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][19][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][20][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][16][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][17][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][18][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][14][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][15][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][16][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][17][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][13][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][14][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][15][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][11][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][12][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][13][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][14][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][10][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][11][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][12][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][8][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][9][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][10][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][11][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][7][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][8][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][9][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[30] <= accum_o_c_30 + accum_o_s_30;

// Coef 31
logic [21:0] accum_i_31 [33];
logic [21:0] accum_o_c_31, accum_o_s_31;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(33),
  .BIT_LEN(22)
)
ct_31 (
  .terms(accum_i_31),
  .C(accum_o_c_31),
  .S(accum_o_s_31)
);
always_comb accum_i_31 = {{{0{1'd0}},mul_grid[5][21][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[5][22][23+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][20][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][21][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[6][22][0+:14],{3{1'd0}}},{{0{1'd0}},mul_grid[7][18][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][19][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][20][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][21][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][17][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][18][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][19][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][15][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][16][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][17][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][18][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][14][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][15][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][16][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][12][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][13][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][14][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][15][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][11][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][12][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][13][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][9][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][10][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][11][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][12][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][8][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][9][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][10][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[31] <= accum_o_c_31 + accum_o_s_31;

// Coef 32
logic [21:0] accum_i_32 [31];
logic [21:0] accum_o_c_32, accum_o_s_32;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(31),
  .BIT_LEN(22)
)
ct_32 (
  .terms(accum_i_32),
  .C(accum_o_c_32),
  .S(accum_o_s_32)
);
always_comb accum_i_32 = {{{0{1'd0}},mul_grid[5][22][40+:3],{0{1'd0}}},{{0{1'd0}},mul_grid[6][21][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[6][22][14+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][19][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][20][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][21][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][22][0+:5],{12{1'd0}}},{{0{1'd0}},mul_grid[8][18][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][19][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][20][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][16][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][17][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][18][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][19][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][15][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][16][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][17][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][13][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][14][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][15][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][16][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][12][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][13][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][14][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][10][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][11][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][12][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][13][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][9][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][10][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][11][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[32] <= accum_o_c_32 + accum_o_s_32;

// Coef 33
logic [21:0] accum_i_33 [28];
logic [21:0] accum_o_c_33, accum_o_s_33;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(28),
  .BIT_LEN(22)
)
ct_33 (
  .terms(accum_i_33),
  .C(accum_o_c_33),
  .S(accum_o_s_33)
);
always_comb accum_i_33 = {{{0{1'd0}},mul_grid[6][22][31+:12],{0{1'd0}}},{{0{1'd0}},mul_grid[7][20][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][21][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[7][22][5+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][19][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][20][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][21][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][17][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][18][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][19][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][20][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][16][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][17][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][18][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][14][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][15][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][16][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][17][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][13][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][14][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][15][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][11][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][12][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][13][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][14][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][10][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][11][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][12][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[33] <= accum_o_c_33 + accum_o_s_33;

// Coef 34
logic [21:0] accum_i_34 [26];
logic [21:0] accum_o_c_34, accum_o_s_34;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(26),
  .BIT_LEN(22)
)
ct_34 (
  .terms(accum_i_34),
  .C(accum_o_c_34),
  .S(accum_o_s_34)
);
always_comb accum_i_34 = {{{0{1'd0}},mul_grid[7][21][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[7][22][22+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][20][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][21][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[8][22][0+:13],{4{1'd0}}},{{0{1'd0}},mul_grid[9][18][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][19][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][20][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][21][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][17][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][18][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][19][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][15][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][16][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][17][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][18][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][14][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][15][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][16][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][12][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][13][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][14][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][15][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][11][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][12][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][13][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[34] <= accum_o_c_34 + accum_o_s_34;

// Coef 35
logic [21:0] accum_i_35 [24];
logic [21:0] accum_o_c_35, accum_o_s_35;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(24),
  .BIT_LEN(22)
)
ct_35 (
  .terms(accum_i_35),
  .C(accum_o_c_35),
  .S(accum_o_s_35)
);
always_comb accum_i_35 = {{{0{1'd0}},mul_grid[7][22][39+:4],{0{1'd0}}},{{0{1'd0}},mul_grid[8][21][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[8][22][13+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][19][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][20][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][21][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][22][0+:4],{13{1'd0}}},{{0{1'd0}},mul_grid[10][18][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][19][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][20][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][16][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][17][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][18][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][19][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][15][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][16][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][17][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][13][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][14][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][15][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][16][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][12][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][13][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][14][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[35] <= accum_o_c_35 + accum_o_s_35;

// Coef 36
logic [21:0] accum_i_36 [21];
logic [21:0] accum_o_c_36, accum_o_s_36;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(21),
  .BIT_LEN(22)
)
ct_36 (
  .terms(accum_i_36),
  .C(accum_o_c_36),
  .S(accum_o_s_36)
);
always_comb accum_i_36 = {{{0{1'd0}},mul_grid[8][22][30+:13],{0{1'd0}}},{{0{1'd0}},mul_grid[9][20][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][21][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[9][22][4+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][19][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][20][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][21][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][17][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][18][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][19][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][20][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][16][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][17][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][18][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][14][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][15][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][16][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][17][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][13][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][14][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][15][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[36] <= accum_o_c_36 + accum_o_s_36;

// Coef 37
logic [20:0] accum_i_37 [19];
logic [20:0] accum_o_c_37, accum_o_s_37;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(19),
  .BIT_LEN(21)
)
ct_37 (
  .terms(accum_i_37),
  .C(accum_o_c_37),
  .S(accum_o_s_37)
);
always_comb accum_i_37 = {{{0{1'd0}},mul_grid[9][21][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[9][22][21+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][20][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][21][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[10][22][0+:12],{5{1'd0}}},{{0{1'd0}},mul_grid[11][18][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][19][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][20][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][21][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][17][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][18][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][19][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][15][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][16][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][17][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][18][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][14][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][15][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][16][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[37] <= accum_o_c_37 + accum_o_s_37;

// Coef 38
logic [20:0] accum_i_38 [17];
logic [20:0] accum_o_c_38, accum_o_s_38;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(17),
  .BIT_LEN(21)
)
ct_38 (
  .terms(accum_i_38),
  .C(accum_o_c_38),
  .S(accum_o_s_38)
);
always_comb accum_i_38 = {{{0{1'd0}},mul_grid[9][22][38+:5],{0{1'd0}}},{{0{1'd0}},mul_grid[10][21][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[10][22][12+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][19][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][20][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][21][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][22][0+:3],{14{1'd0}}},{{0{1'd0}},mul_grid[12][18][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][19][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][20][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][16][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][17][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][18][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][19][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][15][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][16][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][17][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[38] <= accum_o_c_38 + accum_o_s_38;

// Coef 39
logic [20:0] accum_i_39 [14];
logic [20:0] accum_o_c_39, accum_o_s_39;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(14),
  .BIT_LEN(21)
)
ct_39 (
  .terms(accum_i_39),
  .C(accum_o_c_39),
  .S(accum_o_s_39)
);
always_comb accum_i_39 = {{{0{1'd0}},mul_grid[10][22][29+:14],{0{1'd0}}},{{0{1'd0}},mul_grid[11][20][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][21][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[11][22][3+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][19][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][20][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][21][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][17][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][18][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][19][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][20][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][16][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][17][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][18][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[39] <= accum_o_c_39 + accum_o_s_39;

// Coef 40
logic [20:0] accum_i_40 [12];
logic [20:0] accum_o_c_40, accum_o_s_40;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(12),
  .BIT_LEN(21)
)
ct_40 (
  .terms(accum_i_40),
  .C(accum_o_c_40),
  .S(accum_o_s_40)
);
always_comb accum_i_40 = {{{0{1'd0}},mul_grid[11][21][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[11][22][20+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][20][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][21][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[12][22][0+:11],{6{1'd0}}},{{0{1'd0}},mul_grid[13][18][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][19][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][20][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][21][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][17][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][18][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][19][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[40] <= accum_o_c_40 + accum_o_s_40;

// Coef 41
logic [19:0] accum_i_41 [10];
logic [19:0] accum_o_c_41, accum_o_s_41;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(10),
  .BIT_LEN(20)
)
ct_41 (
  .terms(accum_i_41),
  .C(accum_o_c_41),
  .S(accum_o_s_41)
);
always_comb accum_i_41 = {{{0{1'd0}},mul_grid[11][22][37+:6],{0{1'd0}}},{{0{1'd0}},mul_grid[12][21][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[12][22][11+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][19][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][20][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][21][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][22][0+:2],{15{1'd0}}},{{0{1'd0}},mul_grid[14][18][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][19][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][20][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[41] <= accum_o_c_41 + accum_o_s_41;

// Coef 42
logic [19:0] accum_i_42 [7];
logic [19:0] accum_o_c_42, accum_o_s_42;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(7),
  .BIT_LEN(20)
)
ct_42 (
  .terms(accum_i_42),
  .C(accum_o_c_42),
  .S(accum_o_s_42)
);
always_comb accum_i_42 = {{{0{1'd0}},mul_grid[12][22][28+:15],{0{1'd0}}},{{0{1'd0}},mul_grid[13][20][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][21][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[13][22][2+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][19][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][20][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][21][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[42] <= accum_o_c_42 + accum_o_s_42;

// Coef 43
logic [18:0] accum_i_43 [5];
logic [18:0] accum_o_c_43, accum_o_s_43;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(5),
  .BIT_LEN(19)
)
ct_43 (
  .terms(accum_i_43),
  .C(accum_o_c_43),
  .S(accum_o_s_43)
);
always_comb accum_i_43 = {{{0{1'd0}},mul_grid[13][21][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[13][22][19+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][20][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][21][10+:17],{0{1'd0}}},{{0{1'd0}},mul_grid[14][22][0+:10],{7{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[43] <= accum_o_c_43 + accum_o_s_43;

// Coef 44
logic [17:0] accum_i_44 [3];
logic [17:0] accum_o_c_44, accum_o_s_44;
compressor_tree_3_to_2 #(
  .NUM_ELEMENTS(3),
  .BIT_LEN(18)
)
ct_44 (
  .terms(accum_i_44),
  .C(accum_o_c_44),
  .S(accum_o_s_44)
);
always_comb accum_i_44 = {{{0{1'd0}},mul_grid[13][22][36+:7],{0{1'd0}}},{{0{1'd0}},mul_grid[14][21][27+:16],{0{1'd0}}},{{0{1'd0}},mul_grid[14][22][10+:17],{0{1'd0}}}};
always_ff @ (posedge i_clk) accum_grid_o[44] <= accum_o_c_44 + accum_o_s_44;

// Coef 45
always_ff @ (posedge i_clk) accum_grid_o[45] <= {{0{1'd0}},mul_grid[14][22][27+:16],{0{1'd0}}};
